nic specjalnego

*vin wej 0 sin 10 1 1.59k
vin wej 0 pulse 0 1 1n 1n 1n 10us 20us  ; f3 = 6.29ms / 3.14ms	 50kHz to 20us / 10us

*PULSE (V1 V2 TD TR TF PW PER) �
*gdzie    V1 � warto�� pocz�tkowa (w Voltach lub Amperach)
*V2 � warto�� impulsu (w Voltach lub Amperach)
*TD � czas op�nienia (w sekundach, warto�� wbudowana 0.0)
*TR � czas narastania (w sekundach, warto�� wbudowana 0.0)
*TF � czas opadania (w sekundach, warto�� wbudowana 0.0)
*PW � szeroko�� impulsu
*PER � okres impulsu

c1 0 wyj 1u ic=2	   : ic to napi�cie pocz�tkowe na kondensatorze
r1 wej wyj 1k

*.ac dec 100 1000 2000
.tran 1u 0.5m 10u 1u
.probe

.end
